//Модуль для постоянной передачи по Юарт пакетов 
//вида 1 старт-бит =0, 8 бит данных, 1 стоп-бит =1
module cycled_uart_transmitter(
	input 	clk, //Тактовый сигнал
	output reg Tx //Информационный выход
);

// Данные. Максимум 255
parameter data = 8'b1010_1010;

// хранилище данных 10 бит.   
reg [9:0] uart_data;

reg [3:0]i= 1'b0; //счетчик битов = 0

always @ (posedge clk) //с каждым тактом
begin

	//Записываем начальное значение регистра
	uart_data[0] <= 0;//1 старт-бит = 0,
	uart_data[8:1] <= data;//8 бит данных,
	uart_data[9] <= 1;//1 стоп-бит = 1
	
	Tx <= uart_data[i]; //отправили 1 бит данных
	i <= i + 1'b1; //перешли к следующему биту данных
	if(i==9) // если все 10 бит отправлены
	   begin
	     i <= 0;  //обнулить счетчик битов
	   end	
end

endmodule